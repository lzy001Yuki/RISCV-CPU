`include"util.v"
module memory(
    input wire clk,
    input wire rdy_in,
    input wire rst_in,

)
endmodule
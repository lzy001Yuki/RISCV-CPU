`include"util.v"
module predictor(
    input wire clk,
    input wire rdy_in,
    input wire rst_in,

)
endmodule
`include"util.v"
module loadStoreBuffer(
    input wire clk,
    input wire rdy_in,
    input wire rst_in,

)
endmodule